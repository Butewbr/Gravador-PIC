library verilog;
use verilog.vl_types.all;
entity picwriter_tb is
end picwriter_tb;
