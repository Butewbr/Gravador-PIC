library verilog;
use verilog.vl_types.all;
entity halfadder_tb is
end halfadder_tb;
